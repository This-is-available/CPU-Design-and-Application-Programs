`timescale 1ns / 1ns

module pwm_wave_generator(
    input wire clk,
    input wire [15:0] freq,
    output reg signed [9:0] wave_out
);

    reg [5:0] i;
    reg signed [7:0] amplitude [0:63];
    reg [15:0] counter = 0;

    initial begin
        amplitude[0] = 0;
        amplitude[1] = 7;
        amplitude[2] = 13;
        amplitude[3] = 19;
        amplitude[4] = 25;
        amplitude[5] = 30;
        amplitude[6] = 35;
        amplitude[7] = 40;
        amplitude[8] = 45;
        amplitude[9] = 49;
        amplitude[10] = 52;
        amplitude[11] = 55;
        amplitude[12] = 58;
        amplitude[13] = 60;
        amplitude[14] = 62;
        amplitude[15] = 63;
        amplitude[16] = 63;
        amplitude[17] = 63;
        amplitude[18] = 62;
        amplitude[19] = 60;
        amplitude[20] = 58;
        amplitude[21] = 55;
        amplitude[22] = 52;
        amplitude[23] = 49;
        amplitude[24] = 45;
        amplitude[25] = 40;
        amplitude[26] = 35;
        amplitude[27] = 30;
        amplitude[28] = 25;
        amplitude[29] = 19;
        amplitude[30] = 13;
        amplitude[31] = 7;
        amplitude[32] = 0;
        amplitude[33] = -7;
        amplitude[34] = -13;
        amplitude[35] = -19;
        amplitude[36] = -25;
        amplitude[37] = -30;
        amplitude[38] = -35;
        amplitude[39] = -40;
        amplitude[40] = -45;
        amplitude[41] = -49;
        amplitude[42] = -52;
        amplitude[43] = -55;
        amplitude[44] = -58;
        amplitude[45] = -60;
        amplitude[46] = -62;
        amplitude[47] = -63;
        amplitude[48] = -63;
        amplitude[49] = -63;
        amplitude[50] = -62;
        amplitude[51] = -60;
        amplitude[52] = -58;
        amplitude[53] = -55;
        amplitude[54] = -52;
        amplitude[55] = -49;
        amplitude[56] = -45;
        amplitude[57] = -40;
        amplitude[58] = -35;
        amplitude[59] = -30;
        amplitude[60] = -25;
        amplitude[61] = -19;
        amplitude[62] = -13;
        amplitude[63] = -7;
    end

    always @ (posedge clk) begin
      if (freq == 0) wave_out <= 0;
      else if (counter == freq) begin
        counter <= 0;
        wave_out <= $signed(amplitude[i]);
        i <= i + 1;
        if (i == 63) i <= 0; 
        else i <= i + 1;
      end 
      else counter <= counter + 1;
    end
endmodule

module audio_output(
  input wire clk,
  output reg out
);
    wire signed [9:0] ch[0:4];
    wire signed [11:0] wave_sum;
    wire [11:0] positive_wave_sum;
    wire [15:0] freq_count [0:4];
    reg [9:0] PWM;
    reg [31:0] sound [0:79];
    reg [31:0] sound2 [0:79];
    reg [31:0] sound3 [0:180];
    reg [31:0] play_counter;
    reg [15:0] note_counter = 0;
    reg [15:0] note_counter1 = 0;
    reg [31:0] note_data[0:1];
    reg [31:0] note_data2;
    pwm_wave_generator ch0(clk, freq_count[0], ch[0]);
    pwm_wave_generator ch1(clk, freq_count[1], ch[1]);
    pwm_wave_generator ch2(clk, freq_count[2], ch[2]);
    assign freq_count[0] = note_data[0][31:16];
    assign freq_count[1] = note_data[1][31:16];
    assign freq_count[2] = note_data2[31:16];
    assign wave_sum = ch[2] + ch[1] + ch[0];
    assign positive_wave_sum = wave_sum * 2 + 512;
    initial begin
    sound[0] = 32'h0000010a;
    sound[1] = 32'h1284010a;
    sound[2] = 32'h1754010a;
    sound[3] = 32'h18b7010a;
    sound[4] = 32'h0ddf010a;
    sound[5] = 32'h0d17010a;
    sound[6] = 32'h14c80085;
    sound[7] = 32'h0c5b0085;
    sound[8] = 32'h14c80085;
    sound[9] = 32'h00000085;
    sound[10] = 32'h0c5b0085;
    sound[11] = 32'h00000085;
    sound[12] = 32'h0c5b0215;
    sound[13] = 32'h0000010a;
    sound[14] = 32'h0f91026e;
    sound[15] = 32'h000000b1;
    sound[16] = 32'h107f026e;
    sound[17] = 32'h000000b1;
    sound[18] = 32'h0f91026e;
    sound[19] = 32'h00000137;
    sound[20] = 32'h00000085;
    sound[21] = 32'h00000085;
    sound[22] = 32'h00000085;
    sound[23] = 32'h00000085;
    sound[24] = 32'h00000085;
    sound[25] = 32'h0f91026e;
    sound[26] = 32'h000000b1;
    sound[27] = 32'h107f0215;
    sound[28] = 32'h08bd010a;
    sound[29] = 32'h0f91026e;
    sound[30] = 32'h0000034c;
    sound[31] = 32'h00000085;
    sound[32] = 32'h117a026e;
    sound[33] = 32'h000000b1;
    sound[34] = 32'h0b02026e;
    sound[35] = 32'h000000b1;
    sound[36] = 32'h117a026e;
    sound[37] = 32'h00000137;
    sound[38] = 32'h00000085;
    sound[39] = 32'h00000085;
    sound[40] = 32'h00000085;
    sound[41] = 32'h00000085;
    sound[42] = 32'h00000085;
    sound[43] = 32'h0a64026e;
    sound[44] = 32'h000000b1;
    sound[45] = 32'h0f910215;
    sound[46] = 32'h0ddf010a;
    sound[47] = 32'h0f91026e;
    sound[48] = 32'h0000034c;
    sound[49] = 32'h00000085;
    sound[50] = 32'h0942026e;
    sound[51] = 32'h000000b1;
    sound[52] = 32'h07c8026e;
    sound[53] = 32'h000000b1;
    sound[54] = 32'h07c8026e;
    sound[55] = 32'h000000b1;
    sound[56] = 32'h0000010a;
    sound[57] = 32'h00000085;
    sound[58] = 32'h0000010a;
    sound[59] = 32'h00000085;
    sound[60] = 32'h08bd026e;
    sound[61] = 32'h000000b1;
    sound[62] = 32'h08bd026e;
    sound[63] = 32'h000000b1;
    sound[64] = 32'h0baa026e;
    sound[65] = 32'h000000b1;
    sound[66] = 32'h0000010a;
    sound[67] = 32'h00000085;
    sound[68] = 32'h0000010a;
    sound[69] = 32'h00000085;
    sound[70] = 32'h0942026e;
    sound[71] = 32'h000000b1;
    sound[72] = 32'h117a010a;
    sound[73] = 32'h0c5b010a;
    sound[74] = 32'h0c5b010a;
    sound[75] = 32'h09420085;
    sound[76] = 32'h0c5b0085;
    sound[77] = 32'h0942018f;
    sound[78] = 32'h117a0085;
    sound[79] = 32'h1284031f;
    sound2[0] = 32'h14c8010a;
    sound2[1] = 32'h1605010a;
    sound2[2] = 32'h107f010a;
    sound2[3] = 32'h0f91010a;
    sound2[4] = 32'h1754010a;
    sound2[5] = 32'h1605010a;
    sound2[6] = 32'h0c5b0085;
    sound2[7] = 32'h14c80085;
    sound2[8] = 32'h0c5b0085;
    sound2[9] = 32'h00000085;
    sound2[10] = 32'h12840085;
    sound2[11] = 32'h00000085;
    sound2[12] = 32'h117a0215;
    sound2[13] = 32'h0f91010a;
    sound2[14] = 32'h0942026e;
    sound2[15] = 32'h000000b1;
    sound2[16] = 32'h09cf026e;
    sound2[17] = 32'h000000b1;
    sound2[18] = 32'h0942026e;
    sound2[19] = 32'h00000137;
    sound2[20] = 32'h0f910085;
    sound2[21] = 32'h0ddf0085;
    sound2[22] = 32'h0c5b0085;
    sound2[23] = 32'h0baa0085;
    sound2[24] = 32'h0a640085;
    sound2[25] = 32'h0942026e;
    sound2[26] = 32'h000000b1;
    sound2[27] = 32'h09cf0215;
    sound2[28] = 32'h0ddf010a;
    sound2[29] = 32'h0942026e;
    sound2[30] = 32'h0000034c;
    sound2[31] = 32'h0f910085;
    sound2[32] = 32'h0a64026e;
    sound2[33] = 32'h000000b1;
    sound2[34] = 32'h1284026e;
    sound2[35] = 32'h000000b1;
    sound2[36] = 32'h0a64026e;
    sound2[37] = 32'h00000137;
    sound2[38] = 32'h0f910085;
    sound2[39] = 32'h0ddf0085;
    sound2[40] = 32'h0c5b0085;
    sound2[41] = 32'h0baa0085;
    sound2[42] = 32'h0b020085;
    sound2[43] = 32'h117a026e;
    sound2[44] = 32'h000000b1;
    sound2[45] = 32'h18b70215;
    sound2[46] = 32'h08bd010a;
    sound2[47] = 32'h0942026e;
    sound2[48] = 32'h0000034c;
    sound2[49] = 32'h0f910085;
    sound2[50] = 32'h07c8026e;
    sound2[51] = 32'h000000b1;
    sound2[52] = 32'h0a64026e;
    sound2[53] = 32'h000000b1;
    sound2[54] = 32'h0b02026e;
    sound2[55] = 32'h000000b1;
    sound2[56] = 32'h07c8010a;
    sound2[57] = 32'h06ef0085;
    sound2[58] = 32'h0000010a;
    sound2[59] = 32'h07c80085;
    sound2[60] = 32'h0a64026e;
    sound2[61] = 32'h000000b1;
    sound2[62] = 32'h0b02026e;
    sound2[63] = 32'h000000b1;
    sound2[64] = 32'h08bd026e;
    sound2[65] = 32'h000000b1;
    sound2[66] = 32'h08bd010a;
    sound2[67] = 32'h07c80085;
    sound2[68] = 32'h0000010a;
    sound2[69] = 32'h08bd0085;
    sound2[70] = 32'h1754026e;
    sound2[71] = 32'h000000b1;
    sound2[72] = 32'h0ddf010a;
    sound2[73] = 32'h0f91010a;
    sound2[74] = 32'h08bd010a;
    sound2[75] = 32'h0c5b0085;
    sound2[76] = 32'h09420085;
    sound2[77] = 32'h0c5b018f;
    sound2[78] = 32'h0c5b0085;
    sound2[79] = 32'h0baa031f;
    sound3[0] = 32'h00000855;
    sound3[1] = 32'h1f230085;
    sound3[2] = 32'h00000085;
    sound3[3] = 32'h1f23031f;
    sound3[4] = 32'h2ea80085;
    sound3[5] = 32'h00000085;
    sound3[6] = 32'h1f230085;
    sound3[7] = 32'h00000085;
    sound3[8] = 32'h17540085;
    sound3[9] = 32'h00000085;
    sound3[10] = 32'h316e0085;
    sound3[11] = 32'h00000085;
    sound3[12] = 32'h1f230085;
    sound3[13] = 32'h00000085;
    sound3[14] = 32'h18b70085;
    sound3[15] = 32'h00000085;
    sound3[16] = 32'h2ea80085;
    sound3[17] = 32'h00000085;
    sound3[18] = 32'h1f230085;
    sound3[19] = 32'h00000085;
    sound3[20] = 32'h17540085;
    sound3[21] = 32'h00000085;
    sound3[22] = 32'h25080085;
    sound3[23] = 32'h00000085;
    sound3[24] = 32'h1f230085;
    sound3[25] = 32'h00000085;
    sound3[26] = 32'h17540085;
    sound3[27] = 32'h00000085;
    sound3[28] = 32'h2ea80085;
    sound3[29] = 32'h00000085;
    sound3[30] = 32'h1f230085;
    sound3[31] = 32'h00000085;
    sound3[32] = 32'h17540085;
    sound3[33] = 32'h00000085;
    sound3[34] = 32'h316e0085;
    sound3[35] = 32'h00000085;
    sound3[36] = 32'h1f230085;
    sound3[37] = 32'h00000085;
    sound3[38] = 32'h18b70085;
    sound3[39] = 32'h00000085;
    sound3[40] = 32'h2ea80085;
    sound3[41] = 32'h00000085;
    sound3[42] = 32'h1f230085;
    sound3[43] = 32'h00000085;
    sound3[44] = 32'h17540085;
    sound3[45] = 32'h00000085;
    sound3[46] = 32'h25080085;
    sound3[47] = 32'h00000085;
    sound3[48] = 32'h1f230085;
    sound3[49] = 32'h00000085;
    sound3[50] = 32'h17540085;
    sound3[51] = 32'h00000085;
    sound3[52] = 32'h29910085;
    sound3[53] = 32'h00000085;
    sound3[54] = 32'h1f230085;
    sound3[55] = 32'h00000085;
    sound3[56] = 32'h18b70085;
    sound3[57] = 32'h00000085;
    sound3[58] = 32'h2c0a0085;
    sound3[59] = 32'h00000085;
    sound3[60] = 32'h20fe0085;
    sound3[61] = 32'h00000085;
    sound3[62] = 32'h1a2f0085;
    sound3[63] = 32'h00000085;
    sound3[64] = 32'h29910085;
    sound3[65] = 32'h00000085;
    sound3[66] = 32'h1f230085;
    sound3[67] = 32'h00000085;
    sound3[68] = 32'h18b70085;
    sound3[69] = 32'h00000085;
    sound3[70] = 32'h316e0085;
    sound3[71] = 32'h00000085;
    sound3[72] = 32'h1f230085;
    sound3[73] = 32'h00000085;
    sound3[74] = 32'h18b70085;
    sound3[75] = 32'h00000085;
    sound3[76] = 32'h29910085;
    sound3[77] = 32'h00000085;
    sound3[78] = 32'h1f230085;
    sound3[79] = 32'h00000085;
    sound3[80] = 32'h18b70085;
    sound3[81] = 32'h00000085;
    sound3[82] = 32'h316e0085;
    sound3[83] = 32'h00000085;
    sound3[84] = 32'h1f230085;
    sound3[85] = 32'h00000085;
    sound3[86] = 32'h18b70085;
    sound3[87] = 32'h00000085;
    sound3[88] = 32'h2ea80085;
    sound3[89] = 32'h00000085;
    sound3[90] = 32'h1f230085;
    sound3[91] = 32'h00000085;
    sound3[92] = 32'h17540085;
    sound3[93] = 32'h00000085;
    sound3[94] = 32'h3e470085;
    sound3[95] = 32'h00000085;
    sound3[96] = 32'h1f230085;
    sound3[97] = 32'h00000085;
    sound3[98] = 32'h17540085;
    sound3[99] = 32'h00000085;
    sound3[100] = 32'h2ea80085;
    sound3[101] = 32'h00000085;
    sound3[102] = 32'h1f230085;
    sound3[103] = 32'h00000085;
    sound3[104] = 32'h12840085;
    sound3[105] = 32'h00000085;
    sound3[106] = 32'h316e0085;
    sound3[107] = 32'h00000085;
    sound3[108] = 32'h1f230085;
    sound3[109] = 32'h00000085;
    sound3[110] = 32'h14c80085;
    sound3[111] = 32'h00000085;
    sound3[112] = 32'h345f0085;
    sound3[113] = 32'h00000085;
    sound3[114] = 32'h1f230085;
    sound3[115] = 32'h00000085;
    sound3[116] = 32'h16050085;
    sound3[117] = 32'h00000085;
    sound3[118] = 32'h2c0a0085;
    sound3[119] = 32'h00000085;
    sound3[120] = 32'h1f230085;
    sound3[121] = 32'h00000085;
    sound3[122] = 32'h12840085;
    sound3[123] = 32'h00000085;
    sound3[124] = 32'h29910085;
    sound3[125] = 32'h00000085;
    sound3[126] = 32'h1bbe0085;
    sound3[127] = 32'h00000085;
    sound3[128] = 32'h117a0085;
    sound3[129] = 32'h00000085;
    sound3[130] = 32'h2c0a0085;
    sound3[131] = 32'h00000085;
    sound3[132] = 32'h1bbe0085;
    sound3[133] = 32'h00000085;
    sound3[134] = 32'h117a0085;
    sound3[135] = 32'h00000085;
    sound3[136] = 32'h2ea80085;
    sound3[137] = 32'h00000085;
    sound3[138] = 32'h1bbe0085;
    sound3[139] = 32'h00000085;
    sound3[140] = 32'h117a0085;
    sound3[141] = 32'h00000085;
    sound3[142] = 32'h316e0085;
    sound3[143] = 32'h00000085;
    sound3[144] = 32'h1f230085;
    sound3[145] = 32'h00000085;
    sound3[146] = 32'h117a0085;
    sound3[147] = 32'h00000085;
    sound3[148] = 32'h2ea80085;
    sound3[149] = 32'h00000085;
    sound3[150] = 32'h1f230085;
    sound3[151] = 32'h00000085;
    sound3[152] = 32'h12840085;
    sound3[153] = 32'h00000085;
    sound3[154] = 32'h3e470085;
    sound3[155] = 32'h00000085;
    sound3[156] = 32'h1f230085;
    sound3[157] = 32'h00000085;
    sound3[158] = 32'h1f230085;
    sound3[159] = 32'h00000085;
    sound3[160] = 32'h22f40085;
    sound3[161] = 32'h22f40085;
    sound3[162] = 32'h22f4018f;
    sound3[163] = 32'h316e0085;
    sound3[164] = 32'h2ea8031f;

    end
        parameter NOTES = 80;
        parameter BASS = 9'd165;
        parameter PLAY_DELAY = 100_000 - 1;
    always @ (posedge clk) begin
         if (play_counter == PLAY_DELAY) begin
           play_counter <= 0; 
           if (note_data2[15:0] == 0) begin
                   if (note_counter1 == BASS | note_counter1 == 0) begin note_counter1 <= 1; 
                      note_data2 <= sound3[0]; 
                      note_counter <= 1;  note_data[0] <= sound[0];  note_data[1] <= sound2[0];
                      end
                   else begin note_counter1 <= note_counter1 + 1;
                      note_data2 <= sound3[note_counter1]; 
                      end
                   end else note_data2[15:0] <= note_data2[15:0] - 1; 
           if (note_data[0][15:0] == 0) begin
               if (note_counter == 0) begin note_counter <= 1;  note_data[0] <= sound[0];  note_data[1] <= sound2[0];end
               else if (note_counter < NOTES) begin note_counter <= note_counter + 1; note_data[0] <= sound[note_counter];  note_data[1] <= sound2[note_counter]; end
           end else note_data[0][15:0] <= note_data[0][15:0] - 1;
           
         end else play_counter <= play_counter + 1; 
        if (PWM < $unsigned(positive_wave_sum)) out <= 1;
        else out <= 0;
        PWM <= PWM + 1;
    end
endmodule
